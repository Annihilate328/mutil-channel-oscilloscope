module Ms9280_drive(
	Clk,
	Reset_n,
	AD_Clk,
	AD_Data
);
	input Clk;
	input Reset_n;
	output [9:0]AD