module FPGA_oscilloscope(

);


endmodule
