module ADC1_drive(
	input Clk,
	input Reset_n,
	input [7:0] AD_Data,
	input [7:0] Trigger,
	input ADC1_bg,
	input rdreq,
	output reg ADC1_end,
	output empty,
	output [7:0] ADC1_F_O_Data
);
	reg wrreq;
	reg sclr;
	wire full;
	
	// 实例化 ADC0_FIFO
	ADC1_FIFO ADC1_FIFO_inst(
		.clock(Clk),
		.data(AD_Data),
		.rdreq(rdreq),
		.sclr(sclr),
		.wrreq(wrreq),
		.empty(empty),
		.full(full),
		.q(ADC1_F_O_Data),
		.usedw()
	);

	reg [13:0] count;
	reg [2:0] state;
	reg Tri;

	always @(posedge Clk or negedge Reset_n) begin
		if (!Reset_n) begin
			count <= 13'd0;
			ADC1_end <= 0;
		end else begin
			if (count <= 5130) begin
				count <= count + 1'd1;
				if (count >8 && count <1033 && Tri == 1) begin
					count <= 13'd1033;
				end
			end else if (full == 1) begin
				ADC1_end <= 1;
			end else if (ADC1_bg == 1 && empty == 1) begin
				count <= 13'd0;
				ADC1_end <= 0;
			end 
		end
	end

	always @(posedge Clk or negedge Reset_n) begin
		if (!Reset_n) begin
			state <= 3'd0;
		end else begin
			if (count < 9)
				state <= 3'd1;
			else if (count > 8 && count < 1033)
				state <= 3'd2;
			else if(ADC1_end ==1)
				state <= 3'd4;
			else if (count > 1032 && count <5132)
				state <= 3'd3;
			else state <= 3'd0;
		end
	end

	always @(posedge Clk or negedge Reset_n) begin
		if (!Reset_n) begin
			sclr <= 1'b0;
			wrreq <= 1'b0;
		end else begin
			case(state)
				3'd1: begin
					sclr <= 1'b1;
					wrreq <= 1'b0;
				end
				3'd2: begin
					sclr <= 1'b0;
					Tri <= 0;
					if (AD_Data > Trigger && AD_Data < (Trigger + 4'd15)) begin
							Tri <= 1;
					end
				end
				3'd3: begin
					wrreq <= 1'b1;
				end
				3'd4: begin
					wrreq <= 1'b0;
				end
				default: begin
					sclr <= 1'b1;
					Tri <= 1'b0;
					wrreq <= 1'b0;
				end
			endcase
		end
	end
endmodule
